////////////////////////////////////////////////////////////////
// This file houses modules for the inner workings of the ROB //

// This ROB will have 32 entries. We can decide to add or      //
// subtract entries as we see fit.                             //
/////////////////////////////////////////////////////////////////

// parameters //
`define ROB_ENTRIES 32
`define ROB_ENTRY_AVAILABLE 1
`define NO_ROB_ENTRY 0



// rob main module //
module rob(clock,reset, output_value, output_reg, rob_full);

   // inputs //
   input wire clock;
   input wire reset;
   input output_value;
   input output_reg;


   // outputs //
   output rob_full;
   output 




endmodule 

