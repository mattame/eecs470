//////////////////////////////////////////////////////////////////////////
//                                                                      //
//   Modulename :  ex_stage.v                                           //
//                                                                      //
//  Description :  instruction execute (EX) stage of the pipeline;      //
//                 given the instruction command code CMD, select the   //
//                 proper input A and B for the ALU, compute the result,// 
//                 and compute the condition for branches, and pass all //
//                 the results down the pipeline. MWB                   // 
//                                                                      //
//                                                                      //
//////////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps

//
// The Multiplier Stage
//
// given the command code CMD and proper operands A and B, compute the
// result of the instruction
//
// This module is 
//


module mult_stage(clock, reset,
                  product_in,  mplier_in,  mcand_in,  start,
                  product_out, mplier_out, mcand_out, done);

  input clock, reset, start;
  input [63:0] product_in, mplier_in, mcand_in;

  output done;
  output [63:0] product_out, mplier_out, mcand_out;

  reg  [63:0] prod_in_reg, partial_prod_reg;
  wire [63:0] partial_product, next_mplier, next_mcand;

  reg [63:0] mplier_out, mcand_out;
  reg done;

  assign product_out = prod_in_reg + partial_prod_reg;

  assign partial_product = mplier_in[15:0] * mcand_in;

  assign next_mplier = {16'b0,mplier_in[63:16]};
  assign next_mcand = {mcand_in[47:0],16'b0};

  always @(posedge clock)
  begin
    prod_in_reg      <= #1 product_in;
    partial_prod_reg <= #1 partial_product;
    mplier_out       <= #1 next_mplier;
    mcand_out        <= #1 next_mcand;
  end

  always @(posedge clock)
  begin
    if(reset)
      done <= #1 1'b0;
    else
      done <= #1 start;
  end

endmodule                                                                                                                                                                

//
// The Multiplier
//
// given the command code CMD and proper operands A and B, compute the
// product of A and B
//
// This module has four stages, propogating a "done" throughout.
// When the third stage outputs "done", it signals a stall command
// which stalls the pipeline behind it and prevents a structural hazard
// at the end of the EX stage.
//


module mult(clock, reset, mplier, mcand, start, product, stall, done);

  input clock, reset, start;
  input [63:0] mcand, mplier;

  output [63:0] product;
  output done, stall;

  wire [63:0] mcand_out, mplier_out;
  wire [(3*64)-1:0] internal_products, internal_mcands, internal_mpliers;
  wire [1:0] internal_dones;

  mult_stage mstage [3:0]
    (.clock(clock),
     .reset(reset),
     .product_in({internal_products,64'h0}),
     .mplier_in({internal_mpliers,mplier}),
     .mcand_in({internal_mcands,mcand}),
     .start({stall,internal_dones,start}),
     .product_out({product,internal_products}),
     .mplier_out({mplier_out,internal_mpliers}),
     .mcand_out({mcand_out,internal_mcands}),
     .done({done,stall,internal_dones})
    );

endmodule

//
// The ALU
//
// given the command code CMD and proper operands A and B, compute the
// result of the instruction
//
// This module is purely combinational
//

module alu(//Inputs
           opa,
           opb,
           func,
           
           // Output
           result
          );

  input  [63:0] opa;
  input  [63:0] opb;
  input   [4:0] func;
  output [63:0] result;

  reg    [63:0] result;

    // This function computes a signed less-than operation
  function signed_lt;
    input [63:0] a, b;
    
    if (a[63] == b[63]) 
      signed_lt = (a < b); // signs match: signed compare same as unsigned
    else
      signed_lt = a[63];   // signs differ: a is smaller if neg, larger if pos
  endfunction

  always @*
  begin
    case (func)
      `ALU_ADDQ:   result = opa + opb;
      `ALU_SUBQ:   result = opa - opb;
      `ALU_AND:    result = opa & opb;
      `ALU_BIC:    result = opa & ~opb;
      `ALU_BIS:    result = opa | opb;
      `ALU_ORNOT:  result = opa | ~opb;
      `ALU_XOR:    result = opa ^ opb;
      `ALU_EQV:    result = opa ^ ~opb;
      `ALU_SRL:    result = opa >> opb[5:0];
      `ALU_SLL:    result = opa << opb[5:0];
      `ALU_SRA:    result = (opa >> opb[5:0]) | ({64{opa[63]}} << (64 -
                             opb[5:0])); // arithmetic from logical shift
      `ALU_MULQ:   result = opa * opb;
      `ALU_CMPULT: result = { 63'd0, (opa < opb) };
      `ALU_CMPEQ:  result = { 63'd0, (opa == opb) };
      `ALU_CMPULE: result = { 63'd0, (opa <= opb) };
      `ALU_CMPLT:  result = { 63'd0, signed_lt(opa, opb) };
      `ALU_CMPLE:  result = { 63'd0, (signed_lt(opa, opb) || (opa == opb)) };
      default:     result = 64'hdeadbeefbaadbeef; // here only to force
                                                  // a combinational solution
                                                  // a casex would be better
    endcase
  end
endmodule // alu

//
// BrCond module
//
// Given the instruction code, compute the proper condition for the
// instruction; for branches this condition will indicate whether the
// target is taken.
//
// This module is purely combinational
//
module brcond(// Inputs
              opa,        // Value to check against condition
              func,       // Specifies which condition to check

              // Output
              cond        // 0/1 condition result (False/True)
             );

  input   [2:0] func;
  input  [63:0] opa;
  output        cond;
  
  reg           cond;

  always @*
  begin
    case (func[1:0]) // 'full-case'  All cases covered, no need for a default
      2'b00: cond = (opa[0] == 0);  // LBC: (lsb(opa) == 0) ?
      2'b01: cond = (opa == 0);     // EQ: (opa == 0) ?
      2'b10: cond = (opa[63] == 1); // LT: (signed(opa) < 0) : check sign bit
      2'b11: cond = (opa[63] == 1) || (opa == 0); // LE: (signed(opa) <= 0)
    endcase
  
     // negate cond if func[2] is set
    if (func[2])
      cond = ~cond;
  end
endmodule // brcond


module ex_stage(// Inputs
                clock,
                reset,
                id_ex_NPC,
                id_ex_IR,
                id_ex_rega,
                id_ex_regb,
                id_ex_opa_select,
                id_ex_opb_select,
                id_ex_alu_func,
                id_ex_cond_branch,
                id_ex_uncond_branch,
                
                // Outputs
                ex_alu_result_out,
                ex_take_branch_out
               );

  input         clock;               // system clock
  input         reset;               // system reset
  input  [63:0] id_ex_NPC;           // incoming instruction PC+4
  input  [31:0] id_ex_IR;            // incoming instruction
  input  [63:0] id_ex_rega;          // register A value from reg file
  input  [63:0] id_ex_regb;          // register B value from reg file
  input   [1:0] id_ex_opa_select;    // opA mux select from decoder
  input   [1:0] id_ex_opb_select;    // opB mux select from decoder
  input   [4:0] id_ex_alu_func;      // ALU function select from decoder
  input         id_ex_cond_branch;   // is this a cond br? from decoder
  input         id_ex_uncond_branch; // is this an uncond br? from decoder

  output [63:0] ex_alu_result_out;   // ALU result
  output        ex_take_branch_out;  // is this a taken branch?

  reg    [63:0] opa_mux_out, opb_mux_out;
  wire          brcond_result;
   
   // set up possible immediates:
   //   mem_disp: sign-extended 16-bit immediate for memory format
   //   br_disp: sign-extended 21-bit immediate * 4 for branch displacement
   //   alu_imm: zero-extended 8-bit immediate for ALU ops
  wire [63:0] mem_disp = { {48{id_ex_IR[15]}}, id_ex_IR[15:0] };
  wire [63:0] br_disp  = { {41{id_ex_IR[20]}}, id_ex_IR[20:0], 2'b00 };
  wire [63:0] alu_imm  = { 56'b0, id_ex_IR[20:13] };
   
   //
   // ALU opA mux
   //
  always @*
  begin
    case (id_ex_opa_select)
      `ALU_OPA_IS_REGA:     opa_mux_out = id_ex_rega;
      `ALU_OPA_IS_MEM_DISP: opa_mux_out = mem_disp;
      `ALU_OPA_IS_NPC:      opa_mux_out = id_ex_NPC;
      `ALU_OPA_IS_NOT3:     opa_mux_out = ~64'h3;
    endcase
  end

   //
   // ALU opB mux
   //
  always @*
  begin
     // Default value, Set only because the case isnt full.  If you see this
     // value on the output of the mux you have an invalid opb_select
    opb_mux_out = 64'hbaadbeefdeadbeef;
    case (id_ex_opb_select)
      `ALU_OPB_IS_REGB:    opb_mux_out = id_ex_regb;
      `ALU_OPB_IS_ALU_IMM: opb_mux_out = alu_imm;
      `ALU_OPB_IS_BR_DISP: opb_mux_out = br_disp;
    endcase 
  end

   //
   // instantiate the ALU
   //
  alu alu_0 (// Inputs
             .opa(opa_mux_out),
             .opb(opb_mux_out),
             .func(id_ex_alu_func),

             // Output
             .result(ex_alu_result_out)
            );
        
    //
    // instantiate the multiplier
    //

  mult mult_0 (// Inputs
               .clock(clock),
               .reset(reset),
               .mplier(opa_mux_out),
               .mcand(opb_mux_out),
               .start(),
           
               // Outputs
               .product(),
               .stall(),
               .done()
              );
   //
   // instantiate the branch condition tester
   //
  brcond brcond (// Inputs
                .opa(id_ex_rega),       // always check regA value
                .func(id_ex_IR[28:26]), // inst bits to determine check

                // Output
                .cond(brcond_result)
               );

   // ultimate "take branch" signal:
   //    unconditional, or conditional and the condition is true
  assign ex_take_branch_out = id_ex_uncond_branch
                          | (id_ex_cond_branch & brcond_result);

endmodule // module ex_stage

