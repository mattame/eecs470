////////////////////////////////////////////////////////////////
// This file houses modules for the inner workings of the ROB //
////////////////////////////////////////////////////////////////

// parameters //
`define RSTAG_NULL    8'hFF
`define ROB_ENTRIES 8'd16
`define ROB_ENTRY_AVAILABLE 1
`define NO_ROB_ENTRY 0
`define SD #1

// rob entry states //
`define ROBE_EMPTY     2'b00
`define ROBE_INUSE     2'b01
`define ROBE_COMPLETE  2'b10
`define ROBE_UNUSED    2'b11


/***
*   Each ROB Entry needs:
*     State
*     Register to be written to
*     Value to be written
***/
module reorder_buffer_entry(

                  //inputs
                  clock, reset, tag_in
                  register_in, 
                  cdb1_value_in, cdb1_tag_in,
                  cdb2_value_in, cdb2_tag_in,

                  //outputs
                  value_out, register_out, state_out
                  );


  /***  inputs  ***/
  input wire        reset;
  input wire        clock;

  input wire  [7:0] tag_in;

  input wire [63:0] cdb1_value_in, cdb2_value_in;
  input wire  [7:0] cdb1_tag_in, cdb2_tag_in;


  /***  internals  ***/
  reg [63:0]  n_value;
  reg  [4:0]  n_register;
  reg  [1:0]  n_state;
  reg  [1:0]  state;


  /***  outputs  ***/
  output reg [63:0] value_out;
  output reg        complete_out;
  output reg  [4:0] register_out;



  // combinational assignments //  
  always @*
  begin

    //determine whether to latch dispatch
    if (write_enable)
    begin
      n_state    = `ROBE_INUSE;
      n_value    = 64'b0;
      n_register = register_in;
    end

    //determine whether to latch complete 
    else if (~write_enable && tag_in == cdb1_tag_in)
    begin 
      n_state    = `ROBE_COMPLETE;
      n_value    = cdb1_value_in;
      n_register = register_out;
    end
    else if (~write_enable && tag_in == cdb2_tag_in)
    begin
      n_state = `ROBE_COMPLETE;
      n_value = cdb2_value_in;
      n_register = register_out;
    end

    //default case
    else
    begin
      n_state = state_out;
      n_value = value_out;
      n_register = register_out;
    end
  end


  // clock synchronous events //
  always@(posedge clock)
  begin
     if (reset)
     begin
        state_out    <= `SD `ROBE_EMPTY
        value_out    <= `SD 64'h0;
        register_out <= `SD `RSTAG_NULL;
     end
     else
     begin
        state_out    <= `SD n_state;
        value_out    <= `SD n_value;
        register_out <= `SD n_register;
     end


endmodule



/////////////////////
// main ROB module //
/////////////////////
// todo: integrate with rob entry module and set correct inputs for latching
// instruction 
// also, forwarding for the case of a full rob and trying to add instructions
// while retiring is not added, probably should be
module reorder_buffer( clock,reset,
      
      inst1_valid_in,
      inst1_dest_reg,

      inst2_valid_in,
      inst2_dest_reg,

      // tags for reading from the rs // 
      inst1_rega_tag_in,
      inst1_regb_tag_in,
      inst2_rega_tag_in,
      inst2_regb_tag_in,

      // cdb inputs //
      cdb1_tag_in,
      cdb1_value_in,
      cdb2_tag_in,
      cdb2_value_in, 

      // outputs //
      inst1_tag_out,
      inst2_tag_out,

      // values out to the rs //
      inst1_rega_value_out,
      inst1_regb_value_out,
      inst2_rega_value_out,
      inst2_regb_value_out,     

      // signals out //
      rob_full
                 );

   // inputs //
   input wire clock;
   input wire reset; 
   input wire inst1_valid_in;
   input wire inst2_valid_in;
   input wire [4:0] inst1_dest_reg;
   input wire [4:0] inst2_dest_reg;
   input wire [7:0] cdb1_tag_in;
   input wire [7:0] cdb2_tag_in;


   // outputs //
   output wire [7:0] inst1_tag_out;
   output wire [7:0] inst2_tag_out;
   output wire rob_full;


   // internal regs/wires //
   wire [1:0] statuses [(`ROB_ENTRIES-1):0];
   wire [7:0] tail_plus_one; 
   wire [7:0] tail_plus_two;
   reg [7:0]   head;
   reg [7:0] n_head;
   reg [7:0]   tail;
   reg [7:0] n_tail;
   reg   rob_empty;
   reg n_rob_empty;


   // regs/wires for talking directly to ther



   // combinational assignments for head/tail plus one and two. accounts //
   // for overflow  //
   assign head_plus_one = (head==(`ROB_ENTRIES-1)) ? 8'd0 : head+8'd1;
   assign head_plus_two = (head==(`ROB_ENTRIES-1)) ? 8'd1 : ( (head==(`ROB_ENTRIES-2)) ? 8'd0 : head+8'd2 );
   assign tail_plus_one = (tail==(`ROB_ENTRIES-1)) ? 8'd0 : tail+8'd1;                                         
   assign tail_plus_two = (tail==(`ROB_ENTRIES-1)) ? 8'd1 : ( (tail==(`ROB_ENTRIES-2)) ? 8'd0 : tail+8'd2 ); 

   // combinational assignments for signals //
   assign rob_full       = (tail_plus_one==head || tail_plus_two==head); 
   assign inst1_retire   =                  (statuses[head         ]==`ROBE_COMPLETE);
   assign inst2_retire   = (inst1_retire && (statuses[head_plus_one]==`ROBE_COMPLETE) );
   assign inst1_dispatch = ( ~rob_full && (inst1_valid || (~inst1_valid && inst2_valid)) ); 
   assign inst2_dispatch = ( ~rob_full && (inst1_valid && inst2_valid) );


   // combinational assignments for next state signals //
   assign n_head = ( inst1_retire   ? (inst2_retire   ? head_plus_two : head_plus_one) : head );   // if retiring one inst, inc by one. if two, inc by two
   assign n_tail = ( inst1_dispatch ? (inst2_dispatch ? tail_plus_two : tail_plus_one) : tail );   // if dispatching one inst, inc by one. if two, inc by two
   assign n_rob_empty = rob_empty ? ~(tail_plus_one!=head) : 1'b0;   // if empty remain empty unless tail plus one != head, otherwise remain not-empty


   // for tag outputs //
   assign inst1_tag_out = (inst1_dispatch ? tail_plus_one : `RSTAG_NULL);
   assign inst2_tag_out = (inst2_dispatch ? tail_plus_two : `RSTAG_NULL);


   // internal modules for ROB entries //
   genvar i;
   generate 
      for (i=0; i<`ROB_ENTRIES; i=i+1)
      begin

      reservation_station_entry entries ( .clock(clock), .reset(reset),
                                       
                    .tag_in(tags_in[i]),
                    .register_in(registers_in[i]),       
               
                    .cdb1_tag_in(cdb1_tag_in), .cdb1_value_in(cdb1_value_in),
                    .cdb2_tag_in(cdb2_tag_in), .cdb2_value_in(cdb2_value_in),

                    .value_out(values_out[i]),
                    .register_out(registers_out[i]),
                    .state_out(states_out[i])

                         );

      end
   endgenerate


   // clock-synchronouse assignments for //
   always@(posedge clock)
   begin
      if (reset)
      begin
         head      <= 8'd0;
         tail      <= 8'd0;
         rob_empty <= 1'b1;
      end
      else
      begin
         head      <= n_head;
         tail      <= n_tail;
         rob_empty <= n_rob_empty;
      end
   end

endmodule


